
`include "control_signals_struct.svh"

module InstructionExecutor (
    input  logic        clk,                        // Clock signal
    input  logic        reset,                      // Active-low reset
    input  logic [63:0] pc_current,                 // Current PC value (64 bits)
    input  logic [63:0] reg_a_contents,
    input  logic [63:0] reg_b_contents,
    input  control_signals_struct control_signals, 
    input logic execute_enable,
    input logic [63:0] register [31:0],

    output logic [63:0] alu_data_out,               // ALU data output
    output logic [63:0] pc_I_offset_out,            // PC value to jump to
    output  control_signals_struct control_signals_out, 
    output logic        execute_done                // Ready signal indicating execute completion
);


    logic [63:0] ecall_alu_data_out; // Temporary storage for ECALL output
    logic [63:0] alu_result;         // Separate signal for ALU result

    alu ALU_unit(
        .instruction(control_signals.instruction),
        .rs1(reg_a_contents),
        .rs2(reg_b_contents),
        .imm(control_signals.imm),
        .shamt(control_signals.shamt),
        // .alu_enable(alu_enable),
        .pc_alu(pc_current),
        .result(alu_result)
    );

    logic localJumpSignal = 0;
    logic signed [63:0] signed_imm;
    logic [11:0] imm_12bit;
    logic [19:0] imm_20bit;

    logic ecall_done;

    logic [2:0] ecall_counter; // Counter for tracking ECALL cycles (3-bit to count up to 4)
    logic ecall_active;        // Flag to indicate if ECALL is currently active


    always_ff @(posedge clk or posedge reset) begin
        if (reset) begin
            ecall_counter <= 0;
            ecall_active <= 0;
            ecall_done <= 0;
        end else if (execute_enable) begin
            if (control_signals.instruction == 8'd57) begin
                if (!ecall_done && !ecall_active) begin
                    do_ecall(register[17], register[10], register[11], register[12], register[13], register[14], register[15], register[16], ecall_alu_data_out);
                    ecall_active <= 1; // Start ECALL
                    ecall_counter <= 1;
                end else if (ecall_active && ecall_counter < 4) begin
                    ecall_counter <= ecall_counter + 1; // Increment counter
                end else begin
                    ecall_done <= 1; // Set ECALL as done
                    ecall_active <= 0;
                end
            end else begin
                ecall_counter <= 0;
                ecall_active <= 0;
                ecall_done <= 0;
            end
        end
    end



    always_comb begin
        if (reset) begin
            // reg_b_data_out = 64'b0;
            alu_data_out = 64'b0;
            pc_I_offset_out = 64'b0;
            execute_done = 0;
            ecall_alu_data_out = 0;
        end else if (execute_enable) begin
            if(control_signals.opcode == 7'b1100011) begin                      // B-Type Branch (Conditional Jump)
                if (alu_data_out == 1) begin  // branch conditions not met 
                    // Extract the lower 12 bits of the immediate
                    imm_12bit = control_signals.imm[11:0];

                    // Sign-extend the 12-bit immediate to 64 bits
                    
                    signed_imm = {{52{imm_12bit[11]}}, imm_12bit};  // imm_12bit[11] is the sign bit

                    // Perform the addi operation to compute the effective address
                    pc_I_offset_out = control_signals.pc + $signed(signed_imm);
                    localJumpSignal = 1;
                end else begin          // not met
                    pc_I_offset_out = 64'b0;
                    localJumpSignal = 0;
                end
            end else if(control_signals.opcode == 7'b1101111) begin            // JAL J-Type Jump (Unconditional Jump)

                imm_20bit = control_signals.imm[19:0];
                signed_imm = {{44{imm_20bit[19]}}, imm_20bit}; 
                pc_I_offset_out = pc_current + $signed(signed_imm);
                localJumpSignal = 1;

            end else if (control_signals.opcode == 7'b1100111) begin           // I-Type JALR (Unconditional Jump with rs1)

                imm_20bit = control_signals.imm[19:0];
                signed_imm = {{44{imm_20bit[19]}}, imm_20bit}; 
                pc_I_offset_out = reg_a_contents + $signed(signed_imm);
                localJumpSignal = 1;
            
            end else begin
                // no branches, just alu which always runs in comb
                pc_I_offset_out = 64'b0;
                localJumpSignal = 0;
            end
            control_signals_out = control_signals;
            control_signals_out.jump_signal = localJumpSignal;

            if (control_signals.instruction == 8'd57) begin
                alu_data_out = ecall_alu_data_out; // Use ECALL output during operation
            end else begin
                alu_data_out = alu_result; // Default to ALU output
            end

            // Set execute_done based on ECALL state
            if (control_signals.instruction == 8'd57) begin
                if (ecall_done) begin
                    execute_done = 1; // ECALL is fully processed
                end else begin
                    execute_done = 0; // Wait for ECALL to complete
                end
            end else begin
                execute_done = 1; // Non-ECALL instructions always finish in one cycle
            end
        end else begin
            // reg_b_data_out = 64'b0;
            // alu_data_out = 64'b0;
            pc_I_offset_out = 64'b0;
            execute_done = 0;
        end
    end

endmodule